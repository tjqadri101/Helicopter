module clockChecker(clock, clkOut);
	input clock;
	output clkOut;
	
	assign clkOut = clock;

endmodule	